
  library ieee; 
  use ieee.std_logic_1164.all; 
  use ieee.std_logic_unsigned.all; 
  use ieee.std_logic_arith.all;




entity DMA_controller is (
  generic ( 
    adress_width = 32;
    data_width   = 32;
    counter      = 
    
  );
